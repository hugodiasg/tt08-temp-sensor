magic
tech sky130A
magscale 1 2
timestamp 1723763153
<< metal1 >>
rect 810 38440 820 38840
rect 1180 38440 1190 38840
rect 17904 38820 18344 38860
rect 17904 38460 17920 38820
rect 18300 38460 18344 38820
rect 17904 37280 18344 38460
rect 16920 33820 17560 33840
rect 16920 33660 16940 33820
rect 17100 33660 17560 33820
rect 16920 33640 17560 33660
rect 16860 33220 17564 33242
rect 16860 33060 16880 33220
rect 17040 33060 17564 33220
rect 16860 33042 17564 33060
rect 27160 30940 30400 31260
rect 16840 25100 17564 25122
rect 16840 24940 16860 25100
rect 17020 24940 17564 25100
rect 16840 24922 17564 24940
rect 16860 24520 17564 24542
rect 16860 24360 16880 24520
rect 17040 24360 17564 24520
rect 16860 24342 17564 24360
rect 16820 24160 17564 24182
rect 16820 24000 16840 24160
rect 17000 24000 17564 24160
rect 16820 23982 17564 24000
rect 210 23720 220 23920
rect 560 23720 570 23920
rect 16860 23900 17564 23922
rect 16860 23722 16880 23900
rect 16870 23680 16880 23722
rect 17040 23722 17564 23900
rect 17040 23680 17050 23722
rect 30080 1000 30400 30940
rect 30080 720 30100 1000
rect 30380 720 30400 1000
<< via1 >>
rect 820 38440 1180 38840
rect 17920 38460 18300 38820
rect 16940 33660 17100 33820
rect 16880 33060 17040 33220
rect 16860 24940 17020 25100
rect 16880 24360 17040 24520
rect 16840 24000 17000 24160
rect 220 23720 560 23920
rect 16880 23680 17040 23900
rect 30100 720 30380 1000
<< metal2 >>
rect 15220 43820 18960 43840
rect 15220 43660 15240 43820
rect 15400 43660 18820 43820
rect 18920 43660 18960 43820
rect 15220 43640 18960 43660
rect 28740 43120 28820 43130
rect 15900 43080 28740 43100
rect 15900 42920 15920 43080
rect 16080 42920 28740 43080
rect 15900 42900 28740 42920
rect 28820 42900 28840 43100
rect 28740 42890 28820 42900
rect 820 38840 18344 38860
rect 1180 38820 18344 38840
rect 1180 38460 17920 38820
rect 18300 38460 18344 38820
rect 1180 38440 18344 38460
rect 820 38420 18344 38440
rect 13760 33820 17120 33840
rect 13760 33660 13780 33820
rect 13940 33660 16940 33820
rect 17100 33660 17120 33820
rect 13760 33640 17120 33660
rect 14420 33220 17060 33242
rect 14420 33060 14440 33220
rect 14600 33060 16880 33220
rect 17040 33060 17060 33220
rect 14420 33042 17060 33060
rect 15900 25100 17040 25122
rect 15900 24940 15920 25100
rect 16080 24940 16860 25100
rect 17020 24940 17040 25100
rect 15900 24922 17040 24940
rect 15720 24520 17060 24542
rect 15720 24360 15740 24520
rect 15900 24360 16880 24520
rect 17040 24360 17060 24520
rect 15720 24342 17060 24360
rect 15220 24160 17020 24182
rect 15220 24000 15240 24160
rect 15400 24000 16840 24160
rect 17000 24000 17020 24160
rect 15220 23982 17020 24000
rect 220 23922 560 23930
rect 220 23920 17060 23922
rect 560 23900 17060 23920
rect 560 23720 16880 23900
rect 220 23680 16880 23720
rect 17040 23680 17060 23900
rect 220 23620 17060 23680
rect 13760 2940 18960 2960
rect 13760 2780 13780 2940
rect 13940 2780 18780 2940
rect 18940 2780 18960 2940
rect 13760 2760 18960 2780
rect 22640 2260 22820 2270
rect 14420 2240 22640 2260
rect 14420 2080 14440 2240
rect 14600 2080 22640 2240
rect 14420 2060 22820 2080
rect 15720 1740 26700 1760
rect 15720 1580 15740 1740
rect 15900 1580 26500 1740
rect 26680 1580 26700 1740
rect 15720 1560 26700 1580
rect 30100 1000 30380 1010
rect 30100 710 30380 720
<< via2 >>
rect 15240 43660 15400 43820
rect 18820 43660 18920 43820
rect 15920 42920 16080 43080
rect 28740 42900 28820 43120
rect 820 38440 1180 38840
rect 13780 33660 13940 33820
rect 14440 33060 14600 33220
rect 15920 24940 16080 25100
rect 15740 24360 15900 24520
rect 15240 24000 15400 24160
rect 220 23720 560 23920
rect 13780 2780 13940 2940
rect 18780 2780 18940 2940
rect 14440 2080 14600 2240
rect 22640 2080 22820 2260
rect 15740 1580 15900 1740
rect 26500 1580 26680 1740
rect 30100 720 30380 1000
<< metal3 >>
rect 15220 43820 15420 43840
rect 15220 43660 15240 43820
rect 15400 43660 15420 43820
rect 810 38840 1190 38845
rect 810 38440 820 38840
rect 1180 38440 1190 38840
rect 810 38435 1190 38440
rect 13760 33820 13960 33840
rect 13760 33660 13780 33820
rect 13940 33660 13960 33820
rect 210 23920 570 23925
rect 210 23720 220 23920
rect 560 23720 570 23920
rect 210 23715 570 23720
rect 13760 2940 13960 33660
rect 13760 2780 13780 2940
rect 13940 2780 13960 2940
rect 13760 2760 13960 2780
rect 14420 33220 14620 33242
rect 14420 33060 14440 33220
rect 14600 33060 14620 33220
rect 14420 2240 14620 33060
rect 15220 24160 15420 43660
rect 18810 43820 18930 43825
rect 18810 43660 18820 43820
rect 18920 43660 18930 43820
rect 18810 43655 18930 43660
rect 28730 43120 28830 43125
rect 15900 43080 16100 43100
rect 15900 42920 15920 43080
rect 16080 42920 16100 43080
rect 15900 25100 16100 42920
rect 28730 42900 28740 43120
rect 28820 42900 28830 43120
rect 28730 42895 28830 42900
rect 15900 24940 15920 25100
rect 16080 24940 16100 25100
rect 15900 24922 16100 24940
rect 15220 24000 15240 24160
rect 15400 24000 15420 24160
rect 15220 23982 15420 24000
rect 15720 24520 15920 24542
rect 15720 24360 15740 24520
rect 15900 24360 15920 24520
rect 14420 2080 14440 2240
rect 14600 2080 14620 2240
rect 14420 2060 14620 2080
rect 15720 1740 15920 24360
rect 18770 2940 18950 2945
rect 18770 2780 18780 2940
rect 18940 2780 18950 2940
rect 18770 2775 18950 2780
rect 22630 2260 22830 2265
rect 22630 2080 22640 2260
rect 22820 2080 22830 2260
rect 22630 2075 22830 2080
rect 15720 1580 15740 1740
rect 15900 1580 15920 1740
rect 15720 1560 15920 1580
rect 26490 1740 26690 1745
rect 26490 1580 26500 1740
rect 26680 1580 26690 1740
rect 26490 1575 26690 1580
rect 30090 1000 30390 1005
rect 30090 720 30100 1000
rect 30380 720 30390 1000
rect 30090 715 30390 720
<< via3 >>
rect 820 38440 1180 38840
rect 220 23720 560 23920
rect 18820 43660 18920 43820
rect 28740 42900 28820 43120
rect 18780 2780 18940 2940
rect 22640 2080 22820 2260
rect 26500 1580 26680 1740
rect 30100 720 30380 1000
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 200 23920 600 44152
rect 200 23720 220 23920
rect 560 23720 600 23920
rect 200 1000 600 23720
rect 800 38840 1200 44152
rect 18830 43821 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 18819 43820 18921 43821
rect 18819 43660 18820 43820
rect 18920 43660 18921 43820
rect 18819 43659 18921 43660
rect 18830 43650 18890 43659
rect 28766 43121 28826 45152
rect 29318 44952 29378 45152
rect 28739 43120 28826 43121
rect 28739 42900 28740 43120
rect 28820 42900 28826 43120
rect 28739 42899 28826 42900
rect 28766 42890 28826 42899
rect 800 38440 820 38840
rect 1180 38440 1200 38840
rect 800 1000 1200 38440
rect 18770 2940 18950 2970
rect 18770 2780 18780 2940
rect 18940 2780 18950 2940
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 2780
rect 22634 2261 22814 2270
rect 22634 2260 22821 2261
rect 22634 2080 22640 2260
rect 22820 2080 22821 2260
rect 22634 2079 22821 2080
rect 22634 0 22814 2079
rect 26499 1740 26681 1741
rect 26499 1710 26500 1740
rect 26498 1580 26500 1710
rect 26680 1580 26681 1740
rect 26498 1579 26681 1580
rect 26498 0 26678 1579
rect 30050 1000 30542 1010
rect 30050 720 30100 1000
rect 30380 720 30542 1000
rect 30050 670 30542 720
rect 30362 0 30542 670
use device_without_rf  device_without_rf_0 /foss/designs/tt08-temp-sensor/mag/device-complete/mag_without_rf
timestamp 1723762448
transform 0 1 19940 -1 0 38200
box -62 -2580 29620 7540
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 1000 600 44152 1 FreeSans 2 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
